 `timescale 1ns/1ns
module TMA(input [1:0] A, B, input ci, output [1:0] S, output co);
	wire [3:0] p;
	assign p = {A,B};
	assign #(110,91) S[0] = (p == 4'b0000) ? ci :
				 (p == 4'b0001) ? ~ci :
				 (p == 4'b0010) ? ci :
				 (p == 4'b0011) ? ~ci :
				 (p == 4'b0100) ? ~ci :
				 (p == 4'b0101) ? ci :
				 (p == 4'b0110) ? ~ci :
				 (p == 4'b0111) ? ci :
				 (p == 4'b1000) ? ci :
				 (p == 4'b1001) ? ~ci :
				 (p == 4'b1010) ? ci :
				 (p == 4'b1011) ? ~ci :
				 (p == 4'b1100) ? ~ci :
				 (p == 4'b1101) ? ci :
				 (p == 4'b1110) ? ~ci :
				 (p == 4'b1111) ? ci : 1'bx;
	
	assign #(110,91) S[1] = (p == 4'b0000) ? 0 :
				 (p == 4'b0001) ? ci :
				 (p == 4'b0010) ? 1 :
				 (p == 4'b0011) ? ~ci :
				 (p == 4'b0100) ? ci :
				 (p == 4'b0101) ? 1 :
				 (p == 4'b0110) ? ~ci :
				 (p == 4'b0111) ? 0 :
				 (p == 4'b1000) ? 1 :
				 (p == 4'b1001) ? ~ci :
				 (p == 4'b1010) ? 0 :
				 (p == 4'b1011) ? ci :
				 (p == 4'b1100) ? ~ci :
				 (p == 4'b1101) ? 0 :
				 (p == 4'b1110) ? ci :
				 (p == 4'b1111) ? 1 : 1'bx;

	assign #(110,91) co = (p == 4'b0000) ? 0 :
				 (p == 4'b0001) ? 0 :
				 (p == 4'b0010) ? 0 :
				 (p == 4'b0011) ? ci :
				 (p == 4'b0100) ? 0 :
				 (p == 4'b0101) ? 0 :
				 (p == 4'b0110) ? ci :
				 (p == 4'b0111) ? 1 :
				 (p == 4'b1000) ? 0 :
				 (p == 4'b1001) ? ci :
				 (p == 4'b1010) ? 1 :
				 (p == 4'b1011) ? 1 :
				 (p == 4'b1100) ? ci :
				 (p == 4'b1101) ? 1 :
				 (p == 4'b1110) ? 1 :
				 (p == 4'b1111) ? 1 : 1'bx;
endmodule